module BaseCutLine(cut_line,x,y,z);

	parameter LongBits_limit = 10               ; // Sum Of The Data Bit

   //==========================================================================================================
	// Define Type
	//==========================================================================================================	
	typedef bit [LongBits_limit-1:0] LongBitSum ; // Make The LongBitSum Type
	
	//==========================================================================================================
	// Value
	//==========================================================================================================
	int i = 0;
	
	//==========================================================================================================
	// PinData
	//==========================================================================================================
	input  LongBitSum cut_line ; // The Cut Line Ctl Data
	input  LongBitSum x        ; // The Input  X Data
	input  LongBitSum y        ; // The Input  Y Data
	output LongBitSum z        ; // The Output Z Data
	
	//==========================================================================================================
	// Alway Comb Event
	//==========================================================================================================
	always@(*) begin
		for (i=0; i<LongBits_limit; i=i+1) begin
			//Let Two FuzzyNumber Do A Get Min To Max Average
			z[i] = ( (!cut_line[i]) & (x[i] & y[i])) | (cut_line[i] & (x[i] | y[i]));
		end
	end
endmodule
